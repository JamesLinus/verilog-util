//-----------------------------------------------------------------------------
// Title         : A generic linear feedback shift register (random generator)
// Project       : Verilog Utilities
//-----------------------------------------------------------------------------
// File          : lfsr.sv
// Author        : Wei Song  <wsong83@gmail.com>
// Created       : 28.08.2015
// Last modified : 28.08.2015
//-----------------------------------------------------------------------------
//------------------------------------------------------------------------------
// Major modification history :
// 28.08.2015 : created
//-----------------------------------------------------------------------------

module lsfr_seed
  #(
    Length = 8                  // the length of the shifter
    )
   (
    input logic clk, rstn,
    input logic update,         // update the shifter result
    output logic [Length-1:0] data, // the randomized data
    input logic [Length-1:0] seed,  // the seed to be used for initialization, default 0
    input logic seed_valid          // reset seed
    );

   // checking parameters
   initial begin
      assert(Length < 169, "Error: Can generate random data only up to 168 bits!");
      assert(Length > 2, "Error: Can generate random data wider than 2 bits!");
   end

   always_ff @(posedge clk or negedge rstn)
     if(!rstn)
       data <= 0;
     else if(seed_valid)
       data <= seed;
     else if(update)
       data <= lsfr_update(data);

   // see XIlinx document xapp052 for more information
   function logic[Length-1:0] automatic lsfr_update (input logic [Length-1:0] data) begin
      int unsigned eqn [5:0];
      case(Length)
        3:   eqn = '{  3,  2,  0,  0,  0,  0};
        4:   eqn = '{  4,  3,  0,  0,  0,  0};
        5:   eqn = '{  5,  3,  0,  0,  0,  0};
        6:   eqn = '{  6,  5,  0,  0,  0,  0};
        7:   eqn = '{  7,  6,  0,  0,  0,  0};
        8:   eqn = '{  8,  6,  5,  4,  0,  0};
        9:   eqn = '{  9,  5,  0,  0,  0,  0};
        10:  eqn = '{ 10,  7,  0,  0,  0,  0};
        11:  eqn = '{ 11,  9,  0,  0,  0,  0};
        12:  eqn = '{ 12,  6,  4,  1,  0,  0};
        13:  eqn = '{ 13,  4,  3,  1,  0,  0};
        14:  eqn = '{ 14,  5,  3,  1,  0,  0};
        15:  eqn = '{ 15, 14,  0,  0,  0,  0};
        16:  eqn = '{ 16, 15, 13,  4,  0,  0};
        17:  eqn = '{ 17, 14,  0,  0,  0,  0};
        18:  eqn = '{ 18, 11,  0,  0,  0,  0};
        19:  eqn = '{ 19,  6,  2,  1,  0,  0};
        20:  eqn = '{ 20, 17,  0,  0,  0,  0};
        21:  eqn = '{ 21, 19,  0,  0,  0,  0};
        22:  eqn = '{ 22, 21,  0,  0,  0,  0};
        23:  eqn = '{ 23, 18,  0,  0,  0,  0};
        24:  eqn = '{ 24, 23, 22, 17,  0,  0};
        25:  eqn = '{ 25, 22,  0,  0,  0,  0};
        26:  eqn = '{ 26,  6,  2,  1,  0,  0};
        27:  eqn = '{ 27,  5,  2,  1,  0,  0};
        28:  eqn = '{ 28, 25,  0,  0,  0,  0};
        29:  eqn = '{ 29, 27,  0,  0,  0,  0};
        30:  eqn = '{ 30,  6,  4,  1,  0,  0};
        31:  eqn = '{ 31, 28,  0,  0,  0,  0};
        32:  eqn = '{ 32, 22,  2,  1,  0,  0};
        33:  eqn = '{ 33, 20,  0,  0,  0,  0};
        34:  eqn = '{ 34, 27,  2,  1,  0,  0};
        35:  eqn = '{ 35, 33,  0,  0,  0,  0};
        36:  eqn = '{ 36, 25,  0,  0,  0,  0};
        37:  eqn = '{ 37, 5,   4,  3,  2,  1};
        38:  eqn = '{ 38, 6,   5,  1,  0,  0};
        39:  eqn = '{ 39, 35,  0,  0,  0,  0};
        40:  eqn = '{ 40, 38, 21, 19,  0,  0};
        41:  eqn = '{ 41, 38,  0,  0,  0,  0};
        42:  eqn = '{ 42, 41, 20, 19,  0,  0};
        43:  eqn = '{ 43, 42, 38, 37,  0,  0};
        44:  eqn = '{ 44, 43, 18, 17,  0,  0};
        45:  eqn = '{ 45, 44, 42, 41,  0,  0};
        46:  eqn = '{ 46, 45, 26, 25,  0,  0};
        47:  eqn = '{ 47, 42,  0,  0,  0,  0};
        48:  eqn = '{ 48, 47, 21, 20,  0,  0};
        49:  eqn = '{ 49, 40,  0,  0,  0,  0};
        50:  eqn = '{ 50, 49, 24, 23,  0,  0};
        51:  eqn = '{ 51, 50, 36, 35,  0,  0};
        52:  eqn = '{ 52, 49,  0,  0,  0,  0};
        53:  eqn = '{ 53, 52, 38, 37,  0,  0};
        54:  eqn = '{ 54, 53, 18, 17,  0,  0};
        55:  eqn = '{ 55, 31,  0,  0,  0,  0};
        56:  eqn = '{ 56, 55, 35, 34,  0,  0};
        57:  eqn = '{ 57, 50,  0,  0,  0,  0};
        58:  eqn = '{ 58, 39,  0,  0,  0,  0};
        59:  eqn = '{ 59, 58, 38, 37,  0,  0};
        60:  eqn = '{ 60, 59,  0,  0,  0,  0};
        61:  eqn = '{ 61, 60, 46, 45,  0,  0};
        62:  eqn = '{ 62, 61,  6,  5,  0,  0};
        63:  eqn = '{ 63, 62,  0,  0,  0,  0};
        64:  eqn = '{ 64, 63, 61, 60,  0,  0};
        65:  eqn = '{ 65, 47,  0,  0,  0,  0};
        66:  eqn = '{ 66, 65, 57, 56,  0,  0};
        67:  eqn = '{ 67, 66, 58, 57,  0,  0};
        68:  eqn = '{ 68, 59,  0,  0,  0,  0};
        69:  eqn = '{ 69, 67, 42, 40,  0,  0};
        70:  eqn = '{ 70, 69, 55, 54,  0,  0};
        71:  eqn = '{ 71, 65,  0,  0,  0,  0};
        72:  eqn = '{ 72, 66, 25, 19,  0,  0};
        73:  eqn = '{ 73, 48,  0,  0,  0,  0};
        74:  eqn = '{ 74, 73, 59, 58,  0,  0};
        75:  eqn = '{ 75, 74, 65, 64,  0,  0};
        76:  eqn = '{ 76, 75, 41, 40,  0,  0};
        77:  eqn = '{ 77, 76, 47, 46,  0,  0};
        78:  eqn = '{ 78, 77, 59, 58,  0,  0};
        79:  eqn = '{ 79, 70,  0,  0,  0,  0};
        80:  eqn = '{ 80, 79, 43, 42,  0,  0};
        81:  eqn = '{ 81, 77,  0,  0,  0,  0};
        82:  eqn = '{ 82, 79, 47, 44,  0,  0};
        83:  eqn = '{ 83, 82, 38, 37,  0,  0};
        84:  eqn = '{ 84, 71,  0,  0,  0,  0};
        85:  eqn = '{ 85, 84, 58, 57,  0,  0};
        86:  eqn = '{ 86, 85, 74, 73,  0,  0};
        87:  eqn = '{ 87, 74,  0,  0,  0,  0};
        88:  eqn = '{ 88, 87, 17, 16,  0,  0};
        89:  eqn = '{ 89, 51,  0,  0,  0,  0};
        90:  eqn = '{ 90, 89, 72, 71,  0,  0};
        91:  eqn = '{ 91, 90,  8,  7,  0,  0};
        92:  eqn = '{ 92, 91, 80, 79,  0,  0};
        93:  eqn = '{ 93, 91,  0,  0,  0,  0};
        94:  eqn = '{ 94, 73,  0,  0,  0,  0};
        95:  eqn = '{ 95, 84,  0,  0,  0,  0};
        96:  eqn = '{ 96, 94, 49, 47,  0,  0};
        97:  eqn = '{ 97, 91,  0,  0,  0,  0};
        98:  eqn = '{ 98, 87,  0,  0,  0,  0};
        99:  eqn = '{ 99, 97, 54, 52,  0,  0};
        100: eqn = '{100, 63,  0,  0,  0,  0};
        101: eqn = '{101,100, 95, 94,  0,  0};
        102: eqn = '{102,101, 36, 35,  0,  0};
        103: eqn = '{103, 94,  0,  0,  0,  0};
        104: eqn = '{104,103, 94, 93,  0,  0};
        105: eqn = '{105, 89,  0,  0,  0,  0};
        106: eqn = '{106, 91,  0,  0,  0,  0};
        107: eqn = '{107,105, 44, 42,  0,  0};
        108: eqn = '{108, 77,  0,  0,  0,  0};
        109: eqn = '{109,108,103,102,  0,  0};
        110: eqn = '{110,109, 98, 97,  0,  0};
        111: eqn = '{111,101,  0,  0,  0,  0};
        112: eqn = '{112,110, 69, 67,  0,  0};
        113: eqn = '{113,104,  0,  0,  0,  0};
        114: eqn = '{114,113, 33, 32,  0,  0};
        115: eqn = '{115,114,101,100,  0,  0};
        116: eqn = '{116,115, 46, 45,  0,  0};
        117: eqn = '{117,115, 99, 97,  0,  0};
        118: eqn = '{118, 85,  0,  0,  0,  0};
        119: eqn = '{119,111,  0,  0,  0,  0};
        120: eqn = '{120,113,  9,  2,  0,  0};
        121: eqn = '{121,103,  0,  0,  0,  0};
        122: eqn = '{122,121, 63, 62,  0,  0};
        123: eqn = '{123,121,  0,  0,  0,  0};
        124: eqn = '{124, 87,  0,  0,  0,  0};
        125: eqn = '{125,124, 18, 17,  0,  0};
        126: eqn = '{126,125, 90, 89,  0,  0};
        127: eqn = '{127,126,  0,  0,  0,  0};
        128: eqn = '{128,126,101, 99,  0,  0};
        129: eqn = '{129,124,  0,  0,  0,  0};
        130: eqn = '{130,127,  0,  0,  0,  0};
        131: eqn = '{131,130, 84, 83,  0,  0};
        132: eqn = '{132,103,  0,  0,  0,  0};
        133: eqn = '{133,132, 82, 81,  0,  0};
        134: eqn = '{134, 77,  0,  0,  0,  0};
        135: eqn = '{135,124,  0,  0,  0,  0};
        136: eqn = '{136,135, 11, 10,  0,  0};
        137: eqn = '{137,116,  0,  0,  0,  0};
        138: eqn = '{138,137,131,130,  0,  0};
        139: eqn = '{139,136,134,131,  0,  0};
        140: eqn = '{140,111,  0,  0,  0,  0};
        141: eqn = '{141,140,110,109,  0,  0};
        142: eqn = '{142,121,  0,  0,  0,  0};
        143: eqn = '{143,142,123,122,  0,  0};
        144: eqn = '{144,143, 75, 74,  0,  0};
        145: eqn = '{145, 93,  0,  0,  0,  0};
        146: eqn = '{146,145, 87, 86,  0,  0};
        147: eqn = '{147,146,110,109,  0,  0};
        148: eqn = '{148,121,  0,  0,  0,  0};
        149: eqn = '{149,148, 40, 39,  0,  0};
        150: eqn = '{150, 97,  0,  0,  0,  0};
        151: eqn = '{151,148,  0,  0,  0,  0};
        152: eqn = '{152,151, 87, 86,  0,  0};
        153: eqn = '{153,152,  0,  0,  0,  0};
        154: eqn = '{154,152, 27, 25,  0,  0};
        155: eqn = '{155,154,124,123,  0,  0};
        156: eqn = '{156,155, 41, 40,  0,  0};
        157: eqn = '{157,156,131,130,  0,  0};
        158: eqn = '{158,157,132,131,  0,  0};
        159: eqn = '{159,128,  0,  0,  0,  0};
        160: eqn = '{160,159,142,141,  0,  0};
        161: eqn = '{161,143,  0,  0,  0,  0};
        162: eqn = '{162,161, 75, 74,  0,  0};
        163: eqn = '{163,162,104,103,  0,  0};
        164: eqn = '{164,163,151,150,  0,  0};
        165: eqn = '{165,164,135,134,  0,  0};
        166: eqn = '{166,165,128,127,  0,  0};
        167: eqn = '{167,161,  0,  0,  0,  0};
        168: eqn = '{168,166,153,151,  0,  0};
        default:
             eqn = '{  0,  0,  0,  0,  0,  0};
      endcase // case (Length)

      return { data[Length-2],
               eqn[0] == 0 ? 0 : data[Length-eqn[0]] ^
               eqn[1] == 0 ? 0 : data[Length-eqn[1]] ^
               eqn[2] == 0 ? 0 : data[Length-eqn[2]] ^
               eqn[3] == 0 ? 0 : data[Length-eqn[3]] ^
               eqn[4] == 0 ? 0 : data[Length-eqn[4]] ^
               eqn[5] == 0 ? 0 : data[Length-eqn[5]]
               };
   endfunction
 
endmodule // lsfr_seed

// no seed version
module lsfr
  #(
    Length = 8                  // the length of the shifter
    )
   (
    input logic clk, rstn,
    input logic update,         // update the shifter result
    output logic [Length-1:0] data // the randomized data
    );

   lsfr_seed #(Length) U(.*, .seed(0), .seed_valid(1'b0));

endmodule // lsfr
